1,Dutch
2,Other
9,Unknown
