20,"Corop 20"
21,"Corop 21"
21,"Corop 21"
22,"Corop 22"
23,"Corop 23"
24,"Corop 24"
25,"Corop 25"
26,"Corop 26"
27,"Corop 27"
28,"Corop 28"
29,"Corop 29"
30,"Corop 30"
31,"Corop 31"
32,"Corop 32"
33,"Corop 33"
34,"Corop 34"
35,"Corop 35"
36,"Corop 36"
37,"Corop 37"
38,"Corop 38"
38,"Corop 38"
40,"Corop 40"
41,"Corop 41"
 
