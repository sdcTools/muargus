1,male
2,female
