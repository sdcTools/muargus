   1,Aalburg
   2,Aalsmeer
   3,Aalten
   4,Ter Aar
   5,Aardenburg
   6,Aarle-Rixtel
   7,Abcoude
   8,Achtkarspelen
   9,Akersloot
  10,Alblasserdam
  11,Albrandswaard
  12,Alkemade
  13,Alkmaar
  14,Almelo
  15,Almere
  16,Alphen aan den Rijn
  17,Alphen en Riel
  18,Ambt Delden
  19,Ambt Montfort
  20,Ameland
  21,Amerongen
  22,Amersfoort
  23,Ammerzoden
  24,Amstelveen
  25,Amsterdam
  26,Andijk
  27,Angerlo
  28,Anloo
  29,Anna Paulowna
  30,Apeldoorn
  31,Appingedam
  32,Arcen en Velden
  33,Arnemuiden
  34,Arnhem
  35,Assen
  36,Asten
  37,Avereest
  38,Axel
  39,Baarle-Nassau
  40,Baarn
  41,Bakel en Milheeze
  42,Barendrecht
  43,Barneveld
  44,Bathmen
  45,Bedum
  46,Beek
  47,Beek en Donk
  48,Beemster
  49,Beers
  50,Beerta
  51,Beesel
  52,Beilen
  53,Belfeld
  54,Bellingwedde
  55,Bemmel
  56,Bennebroek
  57,Bergambacht
  58,Bergen (L.)
  59,Bergen (NH.)
  60,Bergen op Zoom
  61,Bergeyk
  62,Bergh
  63,Berghem
  64,Bergschenhoek
  65,Berkel en Rodenrijs
  66,Berkel-Enschot
  67,Berlicum
  68,Bernheze@
  69,Bernisse
  70,Best
  71,Beuningen
  72,Beverwijk
  73,het Bildt
  74,Binnenmaas
  75,Bladel en Netersel
  76,Blaricum
  77,Bleiswijk
  78,Bloemendaal
  79,Boarnsterhim
  80,Bodegraven
  81,Boekel
  82,Ten Boer
  83,Bolsward
  84,Borculo
  85,Borger
  86,Born
  87,Borne
  88,Borsele
  89,Boskoop
  90,Boxmeer
  91,Boxtel
  92,Brakel
  93,Breda
  94,Brederwiede
  95,Breukelen
  96,Brielle
  97,Broekhuizen
  98,Brouwershaven
  99,Bruinisse
 100,Brummen
 101,Brunssum
 102,Budel
 103,Bunnik
 104,Bunschoten
 105,Buren
 106,Bussum
 107,Capelle aan den IJssel
 108,Castricum
 109,Chaam
 110,Coevorden
 111,Cothen
 112,Cromstrijen
 113,Cuijk
 114,Cuijk en Sint Agatha
 115,Culemborg
 116,Dalen
 117,Dalfsen
 118,Dantumadeel
 119,De Bilt
 120,De Lier
 121,De Marne
 122,De Ronde Venen
 123,Delft
 124,Delfzijl
 125,Den Dungen
 126,Den Ham
 127,Den Helder
 128,Denekamp
 129,Deurne
 130,Deventer
 131,Didam
 132,Diemen
 133,Diepenheim
 134,Diepenveen
 135,Diessen
 136,Diever
 137,Dinteloord en Prinsenland
 138,Dinxperlo
 139,Dirksland
 140,Dodewaard
 141,Doesburg
 142,Doetinchem
 143,Domburg
 144,Dongen
 145,Dongeradeel
 146,Doorn
 147,Dordrecht
 148,Drechterland
 149,Driebergen-Rijsenburg
 150,Dronten
 151,Drunen
 152,Druten
 153,Duiveland
 154,Duiven
 155,Dussen
 156,Dwingeloo
 157,Echt
 158,Echteld
 159,Edam-Volendam
 160,Ede
 161,Eelde
 162,Eemnes
 163,Eemsmond
 164,Eersel
 165,Egmond
 166,Eibergen
 167,Eijsden
 168,Eindhoven
 169,Elburg
 170,Elst
 171,Emmen
 172,Enkhuizen
 173,Enschede
 174,Epe
 175,Ermelo
 176,Erp
 177,Esch
 178,Etten-Leur
 179,Ferwerderadeel
 180,Fijnaart en Heijningen
 181,Franekeradeel
 182,Gasselte
