1, age under 30
2, age 31-50
3, age 51 and over
8, miss
