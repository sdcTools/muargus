1,Noord
2,Oost
3,West
4,Zuid
