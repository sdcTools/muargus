1,Wheaton
2,Greenham
3,Newbay
4,Oakdale
5,Smokely 
6,Crowdon
7,Mudwater
8,DontKnow
9,Refusal
