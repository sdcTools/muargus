1,Dutch
2,North-Europe
3,South-Europe
4,North-America
5,South-America
6,Mediterrenean
7,African
8,Asian
9,Unknown
