20,Groningen
21,Friesland
22,Drenthe
23,Overijssel
24,Flevoland
25,Gelderland
26,Utrecht
27,Noord-Holland
28,Zuid-Holland
29,Zeeland
30,Noord-Brabant
31,Limburg

