1,regio 1
2,regio 2
3,regio 3
4,regio 4
5,regio 5
6,regio 6
7,regio 7
8,regio 8
9,regio 9
10,regio 10
11,regio 11
12,regio 12
13,regio 13
14,regio 14
15,regio 15
16,regio 16
17,regio 17
18,regio 18

