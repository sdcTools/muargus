1, age under 20
2, age 21-30
3, age 31-40
4, age 41-50
5, age 51-60
6, age 61 and over
